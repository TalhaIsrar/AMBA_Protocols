'timescale 1ns/1ps

module ahb_to_apb_bridge_tb;



endmodule